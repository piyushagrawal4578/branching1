please add verilog code here
